-- control_unit
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity control_unit is
    port(
        clk         : in std_logic;
        rst         : in std_logic;
        opcode      : in std_logic_vector(5 downto 0);   -- op code
        poly_bcd    : in std_logic_vector(15 downto 0);   -- BCD polynomial
        opand1      : in std_logic_vector(15 downto 0);   -- operand 1
        opand2      : in std_logic_vector(15 downto 0);   -- operand 2

        -- registers
        mask        : in  std_logic_vector(15 downto 0);

        -- generation signals
        en_gen      : out std_logic;  -- polynomial generator enable

        -- operation signals
        i           : out std_logic_vector(15 downto 0);  -- i
        j           : out std_logic_vector(15 downto 0);  -- j

        -- memory signals
        mem_data    : in std_logic_vector(15 downto 0);  -- data from memory
        mem_addr    : out std_logic_vector(15 downto 0);  -- address in memory
        mem_t       : inout std_logic;  -- which memory - 0 for elem, 1 for poly
        mem_rd      : out std_logic;  -- read signal to memory

        -- exceptions
        err_b       : out std_logic;  -- out of bound exception
        err_z       : out std_logic  -- zero exception
    );
end control_unit;

architecture structural of control_unit is

    component isbounded
        port(
            operand     : in  std_logic_vector(15 downto 0);
            mask        : in  std_logic_vector(15 downto 0);
            is_out_bd   : out std_logic
        );
    end component;

    component iszero
        port(
            en              : in std_logic;
            operand         : in std_logic_vector(15 downto 0);
            mem_t           : in std_logic;
            is_zero_flag    : out std_logic
        );
    end component;

    signal is_out_bd : std_logic;
    signal en_zero : std_logic;
    signal is_zero_flag : std_logic;
    signal zero_opand : std_logic_vector(15 downto 0);  -- mem_data from memory
    signal bd_opand : std_logic_vector(15 downto 0);  -- mem_data from memory

    type state_type is (op1_state, op2_state);  -- define the states
    signal state : state_type;
    signal temp_data : std_logic_vector(15 downto 0);  -- mem_data from memory

begin

    isbounded_unit: isbounded port map(
        operand => bd_opand,
        mask => mask,
        is_out_bd => err_b
    );

    iszero_unit: iszero port map(
        en => en_zero,
        operand => zero_opand,
        mem_t => mem_t,
        is_zero_flag => err_z
    );

    process (clk, opcode) begin

        if (rising_edge(clk)) then

            case opcode(5 downto 3) is  -- instruction bits

                -- intiate polynomial generator
                when "000" =>

                    -- enable generator
                    en_gen <= '1';

                    -- disable memory lookup
                    mem_t <= 'X';
                    mem_rd <= '0';
                    mem_addr <= "XXXXXXXXXXXXXXXX";

                -- add/sub
                when "001" =>

                    -- disable generator
                    en_gen <= '0';

                    -- disable zero exception
                    en_zero <= '0';

                    case state is

                        when op1_state =>

                            -- if operand 1 is in element form
                            if (opcode(2) = '0') then

                                -- i is converted to polynomial
                                i <= mem_data;

                            -- if operand 1 is in polynomial form
                            else

                                -- i is the user input
                                i <= opand1;
                                bd_opand <= opand1;

                            end if;

                            -- read from memory to convert element to
                            -- polynomial
                            mem_rd <= '1';

                            -- mem2, addr = element, data = polynomial
                            mem_t <= '1';

                            -- address = element
                            mem_addr <= opand2;

                            state <= op2_state;

                        when op2_state =>

                            -- if operand 2 is in element form
                            if (opcode(1) = '0') then

                                -- j is converted to polynomial
                                j <= mem_data;

                            -- if operand 1 is in polynomial form
                            else

                                -- i is the user input
                                j <= opand2;
                                bd_opand <= opand2;

                            end if;

                            state <= op1_state;

                        when others =>

                            -- read from memory to convert element to
                            -- polynomial
                            mem_rd <= '1';

                            -- mem2, addr = element, data = polynomial
                            mem_t <= '1';

                            -- address = element
                            mem_addr <= opand1;

                            -- state initializes to op1_state
                            state <= op1_state;

                    end case;

                -- mul
                when "010" =>

                    -- disable generator
                    en_gen <= '0';

                    -- disable zero exception
                    en_zero <= '0';

                    case state is

                        when op1_state =>

                            -- if operand 1 is in polynomial form
                            if (opcode(2) = '1') then

                                -- i is converted to element
                                i <= mem_data;

                            -- if operand 1 is in element form
                            else

                                -- i is the user input
                                i <= opand1;
                                bd_opand <= opand1;

                            end if;

                            -- read from memory to convert polynomial to
                            -- element
                            mem_rd <= '1';

                            -- mem2, addr = element, data = polynomial
                            mem_t <= '0';

                            -- address = element
                            mem_addr <= opand2;

                            state <= op2_state;

                        when op2_state =>

                            -- if operand 2 is in polynomial form
                            if (opcode(1) = '1') then

                                -- j is converted to element
                                j <= mem_data;

                            -- if operand 1 is in element form
                            else

                                -- i is the user input
                                j <= opand2;
                                bd_opand <= opand2;

                            end if;

                            state <= op1_state;

                        when others =>

                            -- read from memory to convert polynomial to
                            -- element
                            mem_rd <= '1';

                            -- mem1, addr = polynomial, data = element
                            mem_t <= '0';

                            -- address = polynomial
                            mem_addr <= opand1;

                            -- state initializes to op1_state
                            state <= op1_state;

                    end case;

                -- div
                when "011" =>

                    -- disable generator
                    en_gen <= '0';

                    case state is

                        when op1_state =>

                            -- if operand 1 is in polynomial form
                            if (opcode(2) = '1') then

                                -- i is converted to element
                                i <= mem_data;

                            -- if operand 1 is in element form
                            else

                                -- i is the user input
                                i <= opand1;
                                bd_opand <= opand1;

                            end if;

                            -- read from memory to convert polynomial to
                            -- element
                            mem_rd <= '1';

                            -- mem2, addr = element, data = polynomial
                            mem_t <= '0';

                            -- disable zero exception
                            en_zero <= '0';

                            -- address = element
                            mem_addr <= opand2;

                            state <= op2_state;

                        when op2_state =>

                            -- if operand 2 is in polynomial form
                            if (opcode(1) = '1') then

                                -- j is converted to element
                                j <= mem_data;

                                -- disable zero exception
                                en_zero <= '0';

                            -- if operand 1 is in element form
                            else

                                -- i is the user input
                                j <= opand2;
                                bd_opand <= opand2;
                                zero_opand <= opand2;

                                -- enable zero exception
                                en_zero <= '1';

                            end if;

                            state <= op1_state;

                        when others =>

                            -- read from memory to convert polynomial to
                            -- element
                            mem_rd <= '1';

                            -- mem1, addr = polynomial, data = element
                            mem_t <= '0';

                            -- address = polynomial
                            mem_addr <= opand1;

                            -- state initializes to op1_state
                            state <= op1_state;

                    end case;

                -- log
                when "100" =>

                    -- disable generator
                    en_gen <= '0';

                    case state is

                        when op1_state =>

                            -- if operand 1 is in polynomial form
                            if (opcode(2) = '1') then

                                -- i is converted to element
                                i <= mem_data;

                            -- if operand 1 is in element form
                            else

                                -- i is the user input
                                i <= opand1;
                                bd_opand <= opand1;
                                zero_opand <= opand1;

                                -- enable zero exception
                                en_zero <= '1';

                            end if;

                            -- read from memory to convert polynomial to
                            -- element
                            mem_rd <= '1';

                            -- mem2, addr = element, data = polynomial
                            mem_t <= '0';

                            state <= op1_state;

                        when others =>

                            -- read from memory to convert polynomial to
                            -- element
                            mem_rd <= '1';

                            -- mem1, addr = polynomial, data = element
                            mem_t <= '0';

                            -- address = polynomial
                            mem_addr <= opand1;

                            -- state initializes to op1_state
                            state <= op1_state;

                    end case;

                -- reset
                when "101" =>

                    -- disable generator
                    en_gen <= '0';

                    -- disable memory lookup
                    mem_t <= 'X';
                    mem_rd <= '0';
                    mem_addr <= "XXXXXXXXXXXXXXXX";

                -- mode
                when "110" =>

                    -- disable generator
                    en_gen <= '0';

                    -- disable memory lookup
                    mem_t <= 'X';
                    mem_rd <= '0';
                    mem_addr <= "XXXXXXXXXXXXXXXX";

                when "111" =>  -- nop

                    -- disable generator
                    en_gen <= '0';

                    -- disable memory lookup
                    mem_t <= 'X';
                    mem_rd <= '0';
                    mem_addr <= "XXXXXXXXXXXXXXXX";

                when others =>

                    -- disable generator
                    en_gen <= '0';

                    -- disable memory lookup
                    mem_t <= 'X';
                    mem_rd <= '0';
                    mem_addr <= "XXXXXXXXXXXXXXXX";

            end case;

        end if;
        
    end process;

end structural;
